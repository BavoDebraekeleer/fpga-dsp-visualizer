BZh91AY&SY�N: �߀Pyc����������P�qN��\Z ���IOԚa��z����LF&LFA��%%<	��C�4h ��� � ��<yFL��&��d   ��M21M0�&�F	���#C@"�Q<�1&L���x��h��CF�z#�F6$s�ʶ�^'���h����px�?����)X � H .D+
=�$%�H�E�,93����"�k$�t�
::���*wh�_����
F��&�wi���^��K���ٚ.�`�vIQ�k#l{Dr��ʪ[2��W�/����|ubyZ�p�/��Ϗa�D��e2$=�ߕ�Җ!�vu�̡�l�i�8!]�C�ْ1���J��J30�|oT1"�*H�y���iyTܷ�l�#{���0�i��cm�@´�p[���V��V�"�TO	
[%�`���4�X�F+��UFC\����J���:L3�j� ��U������:�� ��>���<�Y���͞%���ۅ��ʍ	0�wY�,�Ɋ�[P�gZH�����4+��ű�[.X1"�
)��ƣv����rJ2/N��s�яp��9��P���ܘ���~��sqK�'q�PMKe¨�{Q	,��L [�vc�P�-��z�XU��a�m���ɤͬh��.�Rؽ�2��v�XN�(ߵ4�Up��0s����z��a��"ʗ���hm���M=�f���Z�8�h<r��8�*m����q�|�~;��Q)�`�!X$�ժ��y1� �A����J!�F�������;�x�>VfpO"[�<��L2d䑍�f����ݳVЕ��]ҁR��X�T�o����$u��u, �X�q@�2��Y�`��yd`�j���`z�5QO�����s�Xa&"H�H�*�b�S�KdL��)B�[��6��xӬ�8�;�HΆ���8k�:3{��|�
�5�J1$����4��4=@�*A�z}Zq��)�s���H�~��F��� �j��\��Ny0�9ݞ�n� ��gPL�@�M�H������W�1���X%��B,]+��z� (�1I�!���\��=� ��n�F�9�J��nv2����a0����|� �i�1�$*���H�
)�'@