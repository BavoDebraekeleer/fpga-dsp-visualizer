BZh91AY&SY^0m` �߀Py����������P����u�	���	���FC@ �  ��&M4�dd�т0�F� H�J��P���i�l����4  @������!� �   $B2L	�����=SM<
hh4z�'�����$�+Ek�'��c��zƉ\BAd_�(!b(����V�vK����!�Nä�QѢ5�c�S�G��D���R0���6��ہ��zR�n�S�Śl��+z��#��0�a$�.��xVm*�o�{��-7�F�a��o�����$$p�*Kr�MصE�-+7%��]���M
Mu!fp�#`�O�{h��w<���3�� 0�F}ł�J�4Χ��n�s-li��cm�@µ(�Ň	�W#Jīqe*'�B��e(��sLE�tf�Z�	�H���H=0"2�`��f��Lc��ֲ�GД������{H̎���؍����="!
���<6k�{,��/b�+�s92Aɳ��ѥ��
G��
!��(�	�d`8Aqp��DM�@���ab/�w$˹��K��[3~��3��~d!xM�d�4�R��	K�@Q\�KYE�'	���%S	F<�T�x��9\9�u-���+�C[�'"(�4�Ul(`��
f����P6�3�R�AY�f��bB!����U��F�۵"�0��7�׸UgHd��������q$��<K��GYP93b$P\�`�ZD���-4V,��������̞2s�W�����YR�3َ��>yT�b�P�(7=ImMD���_0,�
�8�K�bE�0�:LP�J�' D;�e)R�~���34����!��tђ*`R.�#����W��7��>Q���0��*u9�.��p�_z�C���[C5��:���a���,e� nEɗ���MW�:�GB�G���a�XRa`*�����\Rt������e e�۸4�N{�(��T�Q.�Z�BW�Kn�5�b_���q<�p�]�&JU�$�
�&
p���0K����ba-��%�c�r�.�lN�Q%&L��#Sg��Up��A4!�Z�C	�rE8P�^0m`