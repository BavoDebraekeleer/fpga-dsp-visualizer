BZh91AY&SY�^�} �߀Py����߰����P�rJZ�� �QTo�3Q�z���ji�ц��4�!� ��&L��L �0L�0�D)�Lډ���jx��OP4�   ��2b10d�2 h�00	LM6
=M��d�G�2z���IBJ���~��B&�k��y�ўe�jc��&�1��Z��łi4Y��.#V02�ֵ�it�
>�x�FG��I-�⑆�L2p���{R�Q�Pit��"�6���(�!�h�0�H�@!`��U/������~���c�=�l8�Q+��L����hiKBa����TO6.$K��iavk����L��o���̉���XT�����]S>YC�s1���m�q�tY
��0[��<Xv��J��B��eQ��F�
�YU��h����!*4X���Q���1�JU��<�Wu��A�z�g���Nn�(x�@�C��Mi*�!�r6�������nϗ�pa�8���#���kO.�.V�%t���QCF�;4ز6������é�1?h���lDX��Mx#ȑ�tA���g>�Tqa-�s8�@QO��ATR�	�4H�"�ĩӼ�e������=|s-SLJ�@�x�P��4Ye��Rؽ~b��mP�0�F� ���%�At�L�Z���+����+�Cs���/i�l֥a���[5a��+	��&?���.�����=`1s�"8�Ax��C�P�üǁ����$H�P�葴���ݵ\��`�"#yj)�9�(�MA��P𬑡YR�n��hBQ�J� �/��v�e���T���Х�ӤRF6u�
�X
�s��̛���RA�d�I[r���a��<�gt��\�D6��!����h؊�"H��/�ZO���	�؎���B�1Rs5�Er<��]����[Ե�%y�6-	�,M���Cr�.k����f�����V�x����_Xf@�~���qX[`\
��tEA����P�r�\�x��4�5���۸[ǉj��B���Z҅0��ꔴ�da�[t��9�I^a�f���W�H�&�PJ�,���:��d�.=�E��Ԫ��b�vTi�h��a��%�c��bT4���.�p�!��4�